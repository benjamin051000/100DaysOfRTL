module day01 (
	input logic clk, rst,
	input logic d,
	output logic q_no_rst, q_sync_rst, q_async_rst
);

	always_ff @(/* TODO */) begin: dff_no_rst
		
		// TODO your solution here

	end

	always_ff @(/* TODO */) begin: dff_sync_rst

		// TODO your solution here

	end

	always_ff @(/* TODO */) begin: dff_async_rst

		// TODO your solution here
	end

endmodule

