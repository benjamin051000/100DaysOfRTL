 // An edge detector


module day02 (
	input logic clk, rst,
	input logic a,
	output logic rising_edge, falling_edge
);

	// TODO your solution here

endmodule
